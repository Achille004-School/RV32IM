`ifndef RESULT_SRC_VH
`define RESULT_SRC_VH

`define RESULT_SRC_ALU  2'b00
`define RESULT_SRC_LOAD 2'b01
`define RESULT_SRC_PC4  2'b10
`define RESULT_SRC_UNDEFINED 2'bx

`endif