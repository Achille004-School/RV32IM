`ifndef OPCODES_VH
`define OPCODES_VH

// Opcode field values
`define OPCODE_OP      7'b0110011
`define OPCODE_OP_IMM  7'b0010011
`define OPCODE_LOAD    7'b0000011
`define OPCODE_STORE   7'b0100011
`define OPCODE_BRANCH  7'b1100011
`define OPCODE_JALR    7'b1100111
`define OPCODE_JAL     7'b1101111
`define OPCODE_LUI     7'b0110111
`define OPCODE_AUIPC   7'b0010111

`endif